-- spi_pkg.vhd


package spi_pkg is 

	type t_spi_mode is (EXTENDED, DUAL, QUAD);
    type t_dir is (READ, WRITE);

end package;